/*//////////////////////////////////////////////////////////////////////////////////////////////
+--+--+---+-+---+----+
|  |  |   | /   |    |
|  |--|   --    |    |
|  |  |   | \   ---- |
|--+--+---+-+--------+
Module Name:Pkg_64b_Rebuild
Provider:HuKaiLong
Creat Time:2025-03-25 22:46:34
Target Platform:
Function Description: 
//////////////////////////////////////////////////////////////////////////////////////////////*/
`timescale 1ns/1ns


module Pkg_64b_Rebuild (
    input  wire Rst_n,
    input  wire SysClk,

    input  wire logic                    s_clk,
    input  wire logic                    s_rst,

    taxi_axis_if.snk                     s_axis1,
    taxi_axis_if.snk                     s_axis2,

    input  wire logic                    m_clk,
    input  wire logic                    m_rst,
    taxi_axis_if.src                     m_axis


  );
  ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
  ///////////////////////////////////////////            SIGDEF              ////////////////////////////////////////////////////////////
  ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
  // extract parameters
  localparam DATA_W = m_axis.DATA_W;
  localparam logic KEEP_EN = m_axis.KEEP_EN && m_axis.KEEP_EN;
  localparam KEEP_W = m_axis.KEEP_W;
  localparam logic STRB_EN = m_axis.STRB_EN && m_axis.STRB_EN;
  localparam logic LAST_EN = m_axis.LAST_EN && m_axis.LAST_EN;
  localparam logic ID_EN = m_axis.ID_EN && m_axis.ID_EN;
  localparam ID_W = m_axis.ID_W;
  localparam logic DEST_EN = m_axis.DEST_EN && m_axis.DEST_EN;
  localparam DEST_W = m_axis.DEST_W;
  localparam logic USER_EN = m_axis.USER_EN && m_axis.USER_EN;
  localparam USER_W = m_axis.USER_W;

  // check configuration
  if (m_axis.DATA_W != DATA_W)
    $fatal(0, "Error: Interface DATA_W parameter mismatch (instance %m)");

  if (KEEP_EN && m_axis.KEEP_W != KEEP_W)
    $fatal(0, "Error: Interface KEEP_W parameter mismatch (instance %m)");

  ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
  ///////////////////////////////////////////            SUPPORT              ///////////////////////////////////////////////////////////
  ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



  ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
  ///////////////////////////////////////////            LOGIC              /////////////////////////////////////////////////////////////
  ///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



endmodule
